# Swedish translation for bacula-web.
# Copyright (C) 2007 Free Software Foundation, Inc.
# Daniel Nylander <po@danielnylander.se>, 2007.
#
msgid ""
msgstr ""
"Project-Id-Version: bacula-web\n"
"POT-Creation-Date: 2004-06-11 13:02+0200\n"
"PO-Revision-Date: 2007-06-07 17:08+0100\n"
"Last-Translator: Daniel Nylander <po@danielnylander.se>\n"
"Language-Team: Swedish <tp-sv@listor.tp-sv.se>\n"
"MIME-Version: 1.0\n"
"Content-Type: text/plain; charset=utf-8\n"
"Content-Transfer-Encoding: 8bit\n"

#: lang.c:1
#: lang.c:2
msgid "Bytes transferred last 30 days from ALL clients"
msgstr "Byte överförda senaste 30 dagarna från ALLA klienter"

#: lang.c:3
msgid "GENERAL DATA"
msgstr "ALLMÄN DATA"

#: lang.c:4
msgid "Total clients:"
msgstr "Totalt antal klienter:"

#: lang.c:5
msgid "Total bytes stored"
msgstr "Totalt antal byte lagrade"

#: lang.c:6
msgid "Total files:"
msgstr "Totalt antal filer:"

#: lang.c:7
msgid "Last month, bytes transferred"
msgstr "Senast månaden, överförda byte"

#: lang.c:8
msgid "Last month, bytes transferred (pie)"
msgstr "Senast månaden, överförda byte (diagram)"

#: lang.c:9
msgid "General%20report"
msgstr "Allmän%20rapport"

#: lang.c:10
msgid "Status from last 24h"
msgstr "Status senaste 24h"

#: lang.c:11
msgid "Errors:"
msgstr "Fel:"

#: lang.c:12
msgid "Terminated Jobs:"
msgstr "Avbrutna jobb:"

#: lang.c:13
msgid "Total time spent to do backup:"
msgstr "Total tid använd på att göra säkerhetskopior:"

#: lang.c:14
msgid "Bytes transferred last 24h"
msgstr "Byte överförda senaste 24h"

#: lang.c:15
msgid "Show details"
msgstr "Visa detaljer"

#: lang.c:16
msgid "Jobs with errors"
msgstr "Jobb med fel"

#: lang.c:17
msgid "Name"
msgstr "Namn"

#: lang.c:18
msgid "EndTime"
msgstr "Sluttid"

#: lang.c:19
msgid "JobStatus"
msgstr "Jobbstatus"

#: lang.c:20
msgid "Detailed report"
msgstr "Detaljerad rapport"

#: lang.c:21
#: lang.c:42
msgid "Select a job:"
msgstr "Välj ett jobb:"

#: lang.c:22
msgid "go"
msgstr "kör"

#: lang.c:23
msgid "Elapsed time"
msgstr "Återgången tid"

#: lang.c:24
msgid "Job"
msgstr "Jobb"

#: lang.c:25
msgid "Start Time"
msgstr "Starttid"

#: lang.c:26
msgid "End Time"
msgstr "Sluttid"

#: lang.c:27
msgid "Type"
msgstr "Typ"

#: lang.c:28
msgid "Pool"
msgstr "Pool"

#: lang.c:29
#: lang.c:40
msgid "Status"
msgstr "Status"

#: lang.c:30
msgid "Stats Bacula: Job"
msgstr "Statistik Bacula: Jobb"

#: lang.c:31
msgid "Client:"
msgstr "Klient:"

#: lang.c:32
msgid "Period: From"
msgstr "Period: Från"

#: lang.c:33
msgid "to"
msgstr "till"

#: lang.c:34
msgid "Bytes transferred in the period:"
msgstr "Byte överförda under perioden:"

#: lang.c:35
msgid "Files transferred in the period:"
msgstr "Filer överförda under perioden:"

#: lang.c:36
msgid "Date"
msgstr "Datum"

#: lang.c:37
msgid "Elapsed"
msgstr "Återgången"

#: lang.c:38
msgid "Level"
msgstr "Nivå"

#: lang.c:39
msgid "Bytes"
msgstr "Byte"

#: lang.c:41
msgid "SELECT NEW REPORT"
msgstr "VÄLJ NY RAPPORT"

#: lang.c:43
msgid "Graph mode:"
msgstr "Diagramläge:"

#: lang.c:44
msgid "lines"
msgstr "linjer"

#: lang.c:45
msgid "linepoints"
msgstr "linjepunkter"

#: lang.c:46
msgid "points"
msgstr "punkter"

#: lang.c:47
msgid "bars"
msgstr "staplar"

#: lang.c:48
msgid "area"
msgstr "område"

#: lang.c:49
msgid "Data to show:"
msgstr "Data att visa:"

#: lang.c:50
msgid "Transferred bytes"
msgstr "Överförda bytes"

#: lang.c:51
msgid "Start period:"
msgstr "Startperiod:"

#: lang.c:52
msgid "End period:"
msgstr "Slutperiod:"

#: lang.c:53
msgid "Create report"
msgstr "Skapa rapport"

#: lang.c:54
msgid "Volume Name"
msgstr "Volymnamn"

#: lang.c:55
msgid "Volume Bytes"
msgstr "Volymbyte"

#: lang.c:56
msgid "Media Type"
msgstr "Mediatyp"

#: lang.c:57
msgid "When expire?"
msgstr "Förfaller?"

#: lang.c:58
msgid "Last Written"
msgstr "Senast skriven"

#: lang.c:59
msgid "Volume Status"
msgstr "Volymstatus"

